.temp -25.0 0.0 25.0 50.0 75.0 100.0
.param LoadCap = 1f
.param vdd = 0.8
.param number_fin = 5
