.temp -25.0 0.0 25.0 50.0 75.0 100.0 125.0
.param vdd=0.7 
.param vss=0 
.param number_fin = 1
.param LoadCap = 1f
