.temp -25.0
.param load = 1f
.param Vin = 0.9
.param pmosW = 7e-08
.param nmosW = 7e-08
.param passo = 0.01n
.param t_pulse = 2n
.param dl = 0.1p
.param pmosL = 3.2e-08
.param nmosL = 3.2e-08
