.temp -25.0 0.0 25.0 50.0 75.0 100.0
.param vdd=0.7 
.param vss=0 
.param number_fin = 1
.param p_fin = 7*number_fin
.param n_fin = 6*number_fin
.param LoadCap = 1f