.temp -25.0 0.0 25.0 50.0 75.0 100.0 125.0
.param Vin=0.7 
.param vss=0 
.param number_fin = 1
.param load = 1f
.param passo = 0.01n
.param t_pulse = 10n
.param dl = 0.1p
